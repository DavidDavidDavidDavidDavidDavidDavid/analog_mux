magic
tech sky130A
magscale 1 2
timestamp 1683272759
<< nwell >>
rect 5326 749 6141 1070
rect 6698 824 6760 978
rect 5322 -491 5875 -170
rect 6642 -224 6846 -90
rect 6710 -278 6722 -272
rect 6772 -278 6774 -276
rect 6710 -386 6720 -278
rect 6710 -398 6774 -386
rect 5320 -1291 5872 -970
rect 6624 -1018 6856 -906
rect 6662 -1020 6816 -1018
rect 6648 -1820 6856 -1714
rect 6652 -2604 6874 -2500
rect 6652 -3396 6874 -3292
rect 6640 -4222 6862 -4118
rect 6618 -5028 6840 -4924
rect 6622 -5844 6856 -5710
rect 6638 -7006 6860 -6902
<< pwell >>
rect 6484 509 7023 691
rect 6640 424 6848 509
rect 5614 -757 7994 -549
rect 6654 -822 6862 -757
rect 5622 -1557 7908 -1349
rect 6644 -1614 6852 -1557
rect 5470 -2357 7982 -2149
rect 6648 -2422 6856 -2357
rect 5501 -3159 7923 -2949
rect 6640 -3226 6848 -3159
rect 5591 -3963 7925 -3749
rect 6636 -4032 6844 -3963
rect 5550 -4757 7946 -4549
rect 6654 -4818 6862 -4757
rect 5542 -5557 7936 -5349
rect 6648 -5608 6856 -5557
rect 5609 -6367 7873 -6149
rect 6632 -6428 6840 -6367
rect 6507 -7512 6965 -7330
rect 6646 -7594 6854 -7512
<< psubdiff >>
rect 6676 440 6700 474
rect 6750 440 6774 474
rect 6698 -800 6722 -766
rect 6772 -800 6796 -766
rect 6696 -1600 6720 -1566
rect 6770 -1600 6794 -1566
rect 6698 -2400 6722 -2366
rect 6772 -2400 6796 -2366
rect 6698 -3200 6722 -3166
rect 6772 -3200 6796 -3166
rect 6698 -4000 6722 -3966
rect 6772 -4000 6796 -3966
rect 6698 -4800 6722 -4766
rect 6772 -4800 6796 -4766
rect 6698 -5600 6722 -5566
rect 6772 -5600 6796 -5566
rect 6698 -6400 6722 -6366
rect 6772 -6400 6796 -6366
rect 6698 -7582 6722 -7548
rect 6772 -7582 6796 -7548
<< nsubdiff >>
rect 6704 938 6750 962
rect 6704 842 6750 866
rect 6696 -194 6720 -160
rect 6770 -194 6794 -160
rect 6700 -994 6724 -960
rect 6774 -994 6798 -960
rect 6700 -1794 6724 -1760
rect 6774 -1794 6798 -1760
rect 6698 -2592 6722 -2558
rect 6772 -2592 6796 -2558
rect 6698 -3394 6722 -3360
rect 6772 -3394 6796 -3360
rect 6700 -4194 6724 -4160
rect 6774 -4194 6798 -4160
rect 6700 -4994 6724 -4960
rect 6774 -4994 6798 -4960
rect 6698 -5794 6722 -5760
rect 6772 -5794 6796 -5760
rect 6700 -6982 6724 -6948
rect 6774 -6982 6798 -6948
<< psubdiffcont >>
rect 6700 440 6750 474
rect 6722 -800 6772 -766
rect 6720 -1600 6770 -1566
rect 6722 -2400 6772 -2366
rect 6722 -3200 6772 -3166
rect 6722 -4000 6772 -3966
rect 6722 -4800 6772 -4766
rect 6722 -5600 6772 -5566
rect 6722 -6400 6772 -6366
rect 6722 -7582 6772 -7548
<< nsubdiffcont >>
rect 6704 866 6750 938
rect 6720 -194 6770 -160
rect 6724 -994 6774 -960
rect 6724 -1794 6774 -1760
rect 6722 -2592 6772 -2558
rect 6722 -3394 6772 -3360
rect 6724 -4194 6774 -4160
rect 6724 -4994 6774 -4960
rect 6722 -5794 6772 -5760
rect 6724 -6982 6774 -6948
<< locali >>
rect 6565 1015 6815 1049
rect 6704 938 6750 1015
rect 6704 850 6750 866
rect 6565 474 6855 505
rect 6565 471 6700 474
rect 6684 440 6700 471
rect 6750 471 6855 474
rect 6750 440 6766 471
rect 6704 -191 6720 -160
rect 6589 -194 6720 -191
rect 6770 -191 6786 -160
rect 6770 -194 6903 -191
rect 6589 -225 6903 -194
rect 5559 -493 5609 -489
rect 5559 -571 5609 -543
rect 7903 -587 7953 -543
rect 6593 -766 6957 -735
rect 6593 -769 6722 -766
rect 6706 -800 6722 -769
rect 6772 -769 6957 -766
rect 6772 -800 6788 -769
rect 6708 -991 6724 -960
rect 6589 -994 6724 -991
rect 6774 -991 6790 -960
rect 6774 -994 6947 -991
rect 6589 -1025 6947 -994
rect 5560 -1282 5610 -1278
rect 5560 -1360 5610 -1332
rect 7903 -1373 7953 -1327
rect 6595 -1566 6883 -1535
rect 6595 -1569 6720 -1566
rect 6704 -1600 6720 -1569
rect 6770 -1569 6883 -1566
rect 6770 -1600 6786 -1569
rect 6708 -1791 6724 -1760
rect 6589 -1794 6724 -1791
rect 6774 -1791 6790 -1760
rect 6774 -1794 6881 -1791
rect 6589 -1825 6881 -1794
rect 5560 -2082 5610 -2078
rect 5560 -2160 5610 -2132
rect 7903 -2169 7953 -2125
rect 6601 -2366 6911 -2335
rect 6601 -2369 6722 -2366
rect 6706 -2400 6722 -2369
rect 6772 -2369 6911 -2366
rect 6772 -2400 6788 -2369
rect 6706 -2591 6722 -2558
rect 6589 -2592 6722 -2591
rect 6772 -2591 6788 -2558
rect 6772 -2592 6907 -2591
rect 6589 -2625 6907 -2592
rect 5560 -2882 5610 -2878
rect 5560 -2960 5610 -2932
rect 7903 -2971 7953 -2933
rect 6609 -3166 6879 -3135
rect 6609 -3169 6722 -3166
rect 6706 -3200 6722 -3169
rect 6772 -3169 6879 -3166
rect 6772 -3200 6788 -3169
rect 6706 -3391 6722 -3360
rect 6589 -3394 6722 -3391
rect 6772 -3391 6788 -3360
rect 6772 -3394 6923 -3391
rect 6589 -3425 6923 -3394
rect 5560 -3678 5610 -3674
rect 5560 -3756 5610 -3728
rect 7903 -3773 7953 -3731
rect 6595 -3966 6875 -3935
rect 6595 -3969 6722 -3966
rect 6706 -4000 6722 -3969
rect 6772 -3969 6875 -3966
rect 6772 -4000 6788 -3969
rect 6708 -4191 6724 -4160
rect 6589 -4194 6724 -4191
rect 6774 -4191 6790 -4160
rect 6774 -4194 6895 -4191
rect 6589 -4225 6895 -4194
rect 5560 -4474 5610 -4470
rect 5560 -4552 5610 -4524
rect 7903 -4561 7953 -4527
rect 6589 -4766 6889 -4735
rect 6589 -4769 6722 -4766
rect 6706 -4800 6722 -4769
rect 6772 -4769 6889 -4766
rect 6772 -4800 6788 -4769
rect 6708 -4991 6724 -4960
rect 6589 -4994 6724 -4991
rect 6774 -4991 6790 -4960
rect 6774 -4994 6913 -4991
rect 6589 -5025 6913 -4994
rect 5560 -5276 5610 -5272
rect 5560 -5354 5610 -5326
rect 7903 -5369 7953 -5327
rect 6613 -5566 6877 -5535
rect 6613 -5569 6722 -5566
rect 6706 -5600 6722 -5569
rect 6772 -5569 6877 -5566
rect 6772 -5600 6788 -5569
rect 6706 -5791 6722 -5760
rect 6589 -5794 6722 -5791
rect 6772 -5791 6788 -5760
rect 6772 -5794 6891 -5791
rect 6589 -5825 6891 -5794
rect 5560 -6070 5610 -6066
rect 5560 -6148 5610 -6120
rect 7903 -6165 7953 -6137
rect 6535 -6366 6905 -6335
rect 6535 -6369 6722 -6366
rect 6706 -6400 6722 -6369
rect 6772 -6369 6905 -6366
rect 6772 -6400 6788 -6369
rect 6708 -6972 6724 -6948
rect 6593 -6982 6724 -6972
rect 6774 -6972 6790 -6948
rect 6774 -6982 6875 -6972
rect 6593 -7006 6875 -6982
rect 6611 -7548 6843 -7516
rect 6611 -7550 6722 -7548
rect 6706 -7582 6722 -7550
rect 6772 -7550 6843 -7548
rect 6772 -7582 6788 -7550
<< viali >>
rect 5876 754 5946 814
rect 7504 760 7564 820
rect 6046 704 6086 744
rect 6176 704 6216 744
rect 6326 704 6366 744
rect 6456 704 6496 744
rect 6936 704 6976 744
rect 7066 704 7106 744
rect 7216 704 7256 744
rect 7346 704 7386 744
rect 5876 634 5946 694
rect 7503 631 7572 700
rect 5468 -533 5507 -494
rect 5559 -543 5609 -493
rect 7814 -533 7853 -494
rect 7903 -543 7953 -493
rect 5468 -1330 5507 -1291
rect 5560 -1332 5610 -1282
rect 7804 -1333 7843 -1294
rect 7903 -1327 7953 -1277
rect 5466 -2131 5505 -2092
rect 5560 -2132 5610 -2082
rect 7813 -2130 7852 -2091
rect 7903 -2125 7953 -2075
rect 5464 -2931 5503 -2892
rect 5560 -2932 5610 -2882
rect 7808 -2931 7847 -2892
rect 7903 -2933 7953 -2883
rect 5457 -3732 5496 -3693
rect 5560 -3728 5610 -3678
rect 7808 -3733 7847 -3694
rect 7903 -3731 7953 -3681
rect 5466 -4531 5505 -4492
rect 5560 -4524 5610 -4474
rect 7807 -4531 7846 -4492
rect 7903 -4527 7953 -4477
rect 5464 -5330 5503 -5291
rect 5560 -5326 5610 -5276
rect 7802 -5329 7841 -5290
rect 7903 -5327 7953 -5277
rect 5463 -6132 5502 -6093
rect 5560 -6120 5610 -6070
rect 7807 -6134 7846 -6095
rect 7903 -6137 7953 -6087
rect 6634 -7260 6694 -7200
rect 7534 -7260 7594 -7200
rect 6075 -7310 6115 -7270
rect 6205 -7310 6245 -7270
rect 6355 -7310 6395 -7270
rect 6485 -7310 6525 -7270
rect 6963 -7314 7003 -7274
rect 7093 -7314 7133 -7274
rect 7243 -7314 7283 -7274
rect 7373 -7314 7413 -7274
rect 6634 -7388 6694 -7328
rect 7534 -7388 7594 -7328
<< metal1 >>
rect 7700 1080 7900 1168
rect 5036 984 5042 1080
rect 5138 984 7900 1080
rect 7700 968 7900 984
rect 5866 820 5876 824
rect 5864 754 5876 820
rect 5946 820 5956 824
rect 7492 820 7576 826
rect 5946 754 5958 820
rect 7492 760 7504 820
rect 7564 760 7576 820
rect 5864 748 5958 754
rect 6036 754 6096 760
rect 5864 694 5958 700
rect 6034 698 6036 750
rect 6166 754 6226 760
rect 5864 634 5876 694
rect 5946 634 5958 694
rect 6096 698 6098 750
rect 6164 698 6166 750
rect 6316 754 6376 760
rect 6036 688 6096 694
rect 6226 698 6228 750
rect 6314 698 6316 750
rect 6446 754 6506 760
rect 6166 688 6226 694
rect 6376 698 6378 750
rect 6444 698 6446 750
rect 6926 754 6986 760
rect 6316 688 6376 694
rect 6506 698 6508 750
rect 6924 698 6926 750
rect 7056 754 7116 760
rect 6446 688 6506 694
rect 6986 698 6988 750
rect 7054 698 7056 750
rect 7206 754 7266 760
rect 6926 688 6986 694
rect 7116 698 7118 750
rect 7204 698 7206 750
rect 7336 754 7396 760
rect 7492 754 7576 760
rect 7056 688 7116 694
rect 7266 698 7268 750
rect 7334 698 7336 750
rect 7206 688 7266 694
rect 7396 698 7398 750
rect 7491 700 7584 706
rect 7336 688 7396 694
rect 5864 628 5958 634
rect 7491 631 7503 700
rect 7572 631 7584 700
rect 7491 625 7584 631
rect 5500 440 8416 536
rect 8512 440 8518 536
rect 5056 -256 5062 -160
rect 5158 -256 8058 -160
rect 4334 -377 4534 -320
rect 5462 -377 5513 -376
rect 9310 -377 9510 -284
rect 4334 -428 6540 -377
rect 7485 -428 9510 -377
rect 4334 -520 4534 -428
rect 5462 -494 5513 -428
rect 5462 -533 5468 -494
rect 5507 -533 5513 -494
rect 5462 -545 5513 -533
rect 5547 -493 5621 -487
rect 5547 -543 5559 -493
rect 5609 -543 5621 -493
rect 5547 -549 5621 -543
rect 7808 -494 7859 -428
rect 7808 -533 7814 -494
rect 7853 -533 7859 -494
rect 7808 -545 7859 -533
rect 7891 -493 7965 -487
rect 8732 -493 8932 -460
rect 9310 -484 9510 -428
rect 7891 -543 7903 -493
rect 7953 -543 8932 -493
rect 7891 -549 7965 -543
rect 4338 -601 4538 -576
rect 5559 -601 5609 -549
rect 4338 -651 5609 -601
rect 4338 -776 4538 -651
rect 8732 -660 8932 -543
rect 5437 -800 8386 -704
rect 8482 -800 8488 -704
rect 4372 -1177 4572 -1048
rect 5026 -1056 5032 -960
rect 5128 -1056 8058 -960
rect 9206 -1177 9406 -1080
rect 4372 -1228 6540 -1177
rect 7485 -1228 9406 -1177
rect 4372 -1248 4572 -1228
rect 5462 -1291 5513 -1228
rect 5462 -1330 5468 -1291
rect 5507 -1330 5513 -1291
rect 5462 -1342 5513 -1330
rect 5548 -1282 5622 -1276
rect 5548 -1332 5560 -1282
rect 5610 -1332 5622 -1282
rect 5548 -1338 5622 -1332
rect 7798 -1294 7849 -1228
rect 7798 -1333 7804 -1294
rect 7843 -1333 7849 -1294
rect 7891 -1277 7965 -1271
rect 8754 -1277 8954 -1272
rect 7891 -1327 7903 -1277
rect 7953 -1327 8954 -1277
rect 9206 -1280 9406 -1228
rect 7891 -1333 7965 -1327
rect 4376 -1390 4576 -1346
rect 5560 -1390 5610 -1338
rect 7798 -1345 7849 -1333
rect 4376 -1440 5610 -1390
rect 4376 -1546 4576 -1440
rect 8754 -1472 8954 -1327
rect 5436 -1600 8398 -1504
rect 8494 -1600 8500 -1504
rect 5046 -1856 5052 -1760
rect 5148 -1856 8058 -1760
rect 4314 -1977 4514 -1870
rect 9320 -1977 9520 -1892
rect 4314 -2028 6540 -1977
rect 7485 -2028 9520 -1977
rect 4314 -2070 4514 -2028
rect 5460 -2092 5511 -2028
rect 4376 -2190 4576 -2124
rect 5460 -2131 5466 -2092
rect 5505 -2131 5511 -2092
rect 5460 -2143 5511 -2131
rect 5548 -2082 5622 -2076
rect 5548 -2132 5560 -2082
rect 5610 -2132 5622 -2082
rect 5548 -2138 5622 -2132
rect 7807 -2091 7858 -2028
rect 7807 -2130 7813 -2091
rect 7852 -2130 7858 -2091
rect 5560 -2190 5610 -2138
rect 7807 -2142 7858 -2130
rect 7891 -2075 7965 -2069
rect 8814 -2075 9014 -2068
rect 7891 -2125 7903 -2075
rect 7953 -2125 9014 -2075
rect 9320 -2092 9520 -2028
rect 7891 -2131 7965 -2125
rect 4376 -2240 5610 -2190
rect 4376 -2324 4576 -2240
rect 8814 -2268 9014 -2125
rect 5438 -2400 8396 -2304
rect 8492 -2400 8498 -2304
rect 5040 -2655 5046 -2559
rect 5142 -2655 8057 -2559
rect 4336 -2777 4536 -2674
rect 9352 -2777 9552 -2673
rect 4336 -2828 6540 -2777
rect 7485 -2828 9552 -2777
rect 4336 -2876 4536 -2828
rect 5458 -2892 5509 -2828
rect 5458 -2931 5464 -2892
rect 5503 -2931 5509 -2892
rect 5458 -2943 5509 -2931
rect 5548 -2882 5622 -2876
rect 5548 -2932 5560 -2882
rect 5610 -2932 5622 -2882
rect 5548 -2938 5622 -2932
rect 7802 -2892 7853 -2828
rect 9352 -2873 9552 -2828
rect 7802 -2931 7808 -2892
rect 7847 -2931 7853 -2892
rect 4366 -2990 4566 -2948
rect 5560 -2990 5610 -2938
rect 7802 -2943 7853 -2931
rect 7891 -2883 7965 -2877
rect 8842 -2883 9042 -2882
rect 7891 -2933 7903 -2883
rect 7953 -2933 9042 -2883
rect 7891 -2939 7965 -2933
rect 4366 -3040 5610 -2990
rect 4366 -3148 4566 -3040
rect 8842 -3082 9042 -2933
rect 5437 -3200 8380 -3104
rect 8476 -3200 8482 -3104
rect 4356 -3577 4556 -3436
rect 5056 -3456 5062 -3360
rect 5158 -3456 8056 -3360
rect 9320 -3577 9520 -3454
rect 4356 -3628 6540 -3577
rect 7485 -3628 9520 -3577
rect 4356 -3636 4556 -3628
rect 5451 -3693 5502 -3628
rect 4366 -3786 4566 -3696
rect 5451 -3732 5457 -3693
rect 5496 -3732 5502 -3693
rect 5451 -3744 5502 -3732
rect 5548 -3678 5622 -3672
rect 5548 -3728 5560 -3678
rect 5610 -3728 5622 -3678
rect 5548 -3734 5622 -3728
rect 7802 -3694 7853 -3628
rect 9320 -3654 9520 -3628
rect 7802 -3733 7808 -3694
rect 7847 -3733 7853 -3694
rect 5560 -3786 5610 -3734
rect 7802 -3745 7853 -3733
rect 7891 -3681 7965 -3675
rect 8862 -3681 9062 -3664
rect 7891 -3731 7903 -3681
rect 7953 -3731 9062 -3681
rect 7891 -3737 7965 -3731
rect 4366 -3836 5610 -3786
rect 4366 -3896 4566 -3836
rect 8862 -3864 9062 -3731
rect 5436 -4000 8370 -3904
rect 8466 -4000 8472 -3904
rect 5030 -4256 5036 -4160
rect 5132 -4256 8057 -4160
rect 4348 -4377 4548 -4260
rect 9246 -4377 9446 -4270
rect 4348 -4428 6540 -4377
rect 7485 -4428 9446 -4377
rect 4348 -4460 4548 -4428
rect 5460 -4492 5511 -4428
rect 5460 -4531 5466 -4492
rect 5505 -4531 5511 -4492
rect 5548 -4474 5622 -4468
rect 5548 -4524 5560 -4474
rect 5610 -4524 5622 -4474
rect 5548 -4530 5622 -4524
rect 7801 -4492 7852 -4428
rect 5460 -4543 5511 -4531
rect 4386 -4582 4586 -4552
rect 5560 -4582 5610 -4530
rect 7801 -4531 7807 -4492
rect 7846 -4531 7852 -4492
rect 7801 -4543 7852 -4531
rect 7891 -4477 7965 -4471
rect 8878 -4477 9078 -4466
rect 9246 -4470 9446 -4428
rect 7891 -4527 7903 -4477
rect 7953 -4527 9078 -4477
rect 7891 -4533 7965 -4527
rect 4386 -4632 5610 -4582
rect 4386 -4752 4586 -4632
rect 8878 -4666 9078 -4527
rect 5437 -4800 8388 -4704
rect 8484 -4800 8490 -4704
rect 5030 -5056 5036 -4960
rect 5132 -5056 8058 -4960
rect 4350 -5177 4550 -5110
rect 9374 -5177 9574 -5035
rect 4350 -5228 6540 -5177
rect 7485 -5228 9574 -5177
rect 4350 -5310 4550 -5228
rect 5458 -5291 5509 -5228
rect 5458 -5330 5464 -5291
rect 5503 -5330 5509 -5291
rect 5458 -5342 5509 -5330
rect 5548 -5276 5622 -5270
rect 5548 -5326 5560 -5276
rect 5610 -5326 5622 -5276
rect 5548 -5332 5622 -5326
rect 7796 -5290 7847 -5228
rect 9374 -5235 9574 -5228
rect 7796 -5329 7802 -5290
rect 7841 -5329 7847 -5290
rect 4356 -5384 4556 -5358
rect 5560 -5384 5610 -5332
rect 7796 -5341 7847 -5329
rect 7891 -5277 7965 -5271
rect 8942 -5277 9142 -5266
rect 7891 -5327 7903 -5277
rect 7953 -5327 9142 -5277
rect 7891 -5333 7965 -5327
rect 4356 -5434 5610 -5384
rect 4356 -5558 4556 -5434
rect 8942 -5466 9142 -5327
rect 5435 -5600 8370 -5504
rect 8466 -5600 8472 -5504
rect 4324 -5977 4524 -5836
rect 5026 -5856 5032 -5760
rect 5128 -5856 8057 -5760
rect 9354 -5977 9554 -5848
rect 4324 -6028 6540 -5977
rect 7485 -6028 9554 -5977
rect 4324 -6036 4524 -6028
rect 5457 -6093 5508 -6028
rect 4366 -6178 4566 -6124
rect 5457 -6132 5463 -6093
rect 5502 -6132 5508 -6093
rect 5548 -6070 5622 -6064
rect 5548 -6120 5560 -6070
rect 5610 -6120 5622 -6070
rect 5548 -6126 5622 -6120
rect 7801 -6095 7852 -6028
rect 9354 -6048 9554 -6028
rect 5457 -6144 5508 -6132
rect 5560 -6178 5610 -6126
rect 7801 -6134 7807 -6095
rect 7846 -6134 7852 -6095
rect 7801 -6146 7852 -6134
rect 7891 -6087 7965 -6081
rect 8892 -6087 9092 -6060
rect 7891 -6137 7903 -6087
rect 7953 -6137 9092 -6087
rect 7891 -6143 7965 -6137
rect 4366 -6228 5610 -6178
rect 4366 -6324 4566 -6228
rect 8892 -6260 9092 -6137
rect 5437 -6399 8394 -6303
rect 8490 -6399 8496 -6303
rect 5026 -7044 5032 -6948
rect 5128 -7044 7956 -6948
rect 6622 -7200 6706 -7194
rect 6065 -7260 6125 -7254
rect 6063 -7316 6065 -7264
rect 6195 -7260 6255 -7254
rect 6125 -7316 6127 -7264
rect 6193 -7316 6195 -7264
rect 6345 -7260 6405 -7254
rect 6065 -7326 6125 -7320
rect 6255 -7316 6257 -7264
rect 6343 -7316 6345 -7264
rect 6475 -7260 6535 -7254
rect 6195 -7326 6255 -7320
rect 6405 -7316 6407 -7264
rect 6473 -7316 6475 -7264
rect 6622 -7260 6634 -7200
rect 6694 -7260 6706 -7200
rect 7522 -7200 7606 -7194
rect 6345 -7326 6405 -7320
rect 6535 -7316 6537 -7264
rect 6622 -7266 6706 -7260
rect 6953 -7264 7013 -7258
rect 6951 -7320 6953 -7268
rect 7083 -7264 7143 -7258
rect 6475 -7326 6535 -7320
rect 6622 -7328 6706 -7322
rect 6622 -7388 6634 -7328
rect 6694 -7388 6706 -7328
rect 7013 -7320 7015 -7268
rect 7081 -7320 7083 -7268
rect 7233 -7264 7293 -7258
rect 6953 -7330 7013 -7324
rect 7143 -7320 7145 -7268
rect 7231 -7320 7233 -7268
rect 7363 -7264 7423 -7258
rect 7083 -7330 7143 -7324
rect 7293 -7320 7295 -7268
rect 7361 -7320 7363 -7268
rect 7522 -7260 7534 -7200
rect 7594 -7260 7606 -7200
rect 7522 -7266 7606 -7260
rect 7233 -7330 7293 -7324
rect 7423 -7320 7425 -7268
rect 7363 -7330 7423 -7324
rect 7522 -7328 7606 -7322
rect 6622 -7394 6706 -7388
rect 7522 -7388 7534 -7328
rect 7594 -7388 7606 -7328
rect 7522 -7394 7606 -7388
rect 5606 -7486 5806 -7434
rect 5606 -7582 8372 -7486
rect 8468 -7582 8474 -7486
rect 5606 -7634 5806 -7582
<< via1 >>
rect 5042 984 5138 1080
rect 5876 814 5946 824
rect 5876 764 5946 814
rect 7504 760 7564 820
rect 6036 744 6096 754
rect 6036 704 6046 744
rect 6046 704 6086 744
rect 6086 704 6096 744
rect 5876 634 5946 694
rect 6036 694 6096 704
rect 6166 744 6226 754
rect 6166 704 6176 744
rect 6176 704 6216 744
rect 6216 704 6226 744
rect 6166 694 6226 704
rect 6316 744 6376 754
rect 6316 704 6326 744
rect 6326 704 6366 744
rect 6366 704 6376 744
rect 6316 694 6376 704
rect 6446 744 6506 754
rect 6446 704 6456 744
rect 6456 704 6496 744
rect 6496 704 6506 744
rect 6446 694 6506 704
rect 6926 744 6986 754
rect 6926 704 6936 744
rect 6936 704 6976 744
rect 6976 704 6986 744
rect 6926 694 6986 704
rect 7056 744 7116 754
rect 7056 704 7066 744
rect 7066 704 7106 744
rect 7106 704 7116 744
rect 7056 694 7116 704
rect 7206 744 7266 754
rect 7206 704 7216 744
rect 7216 704 7256 744
rect 7256 704 7266 744
rect 7206 694 7266 704
rect 7336 744 7396 754
rect 7336 704 7346 744
rect 7346 704 7386 744
rect 7386 704 7396 744
rect 7336 694 7396 704
rect 7503 631 7572 700
rect 8416 440 8512 536
rect 5062 -256 5158 -160
rect 8386 -800 8482 -704
rect 5032 -1056 5128 -960
rect 8398 -1600 8494 -1504
rect 5052 -1856 5148 -1760
rect 8396 -2400 8492 -2304
rect 5046 -2655 5142 -2559
rect 8380 -3200 8476 -3104
rect 5062 -3456 5158 -3360
rect 8370 -4000 8466 -3904
rect 5036 -4256 5132 -4160
rect 8388 -4800 8484 -4704
rect 5036 -5056 5132 -4960
rect 8370 -5600 8466 -5504
rect 5032 -5856 5128 -5760
rect 8394 -6399 8490 -6303
rect 5032 -7044 5128 -6948
rect 6065 -7270 6125 -7260
rect 6065 -7310 6075 -7270
rect 6075 -7310 6115 -7270
rect 6115 -7310 6125 -7270
rect 6065 -7320 6125 -7310
rect 6195 -7270 6255 -7260
rect 6195 -7310 6205 -7270
rect 6205 -7310 6245 -7270
rect 6245 -7310 6255 -7270
rect 6195 -7320 6255 -7310
rect 6345 -7270 6405 -7260
rect 6345 -7310 6355 -7270
rect 6355 -7310 6395 -7270
rect 6395 -7310 6405 -7270
rect 6345 -7320 6405 -7310
rect 6475 -7270 6535 -7260
rect 6634 -7260 6694 -7200
rect 6475 -7310 6485 -7270
rect 6485 -7310 6525 -7270
rect 6525 -7310 6535 -7270
rect 6475 -7320 6535 -7310
rect 6953 -7274 7013 -7264
rect 6953 -7314 6963 -7274
rect 6963 -7314 7003 -7274
rect 7003 -7314 7013 -7274
rect 6634 -7388 6694 -7328
rect 6953 -7324 7013 -7314
rect 7083 -7274 7143 -7264
rect 7083 -7314 7093 -7274
rect 7093 -7314 7133 -7274
rect 7133 -7314 7143 -7274
rect 7083 -7324 7143 -7314
rect 7233 -7274 7293 -7264
rect 7233 -7314 7243 -7274
rect 7243 -7314 7283 -7274
rect 7283 -7314 7293 -7274
rect 7233 -7324 7293 -7314
rect 7363 -7274 7423 -7264
rect 7534 -7260 7594 -7200
rect 7363 -7314 7373 -7274
rect 7373 -7314 7413 -7274
rect 7413 -7314 7423 -7274
rect 7363 -7324 7423 -7314
rect 7534 -7388 7594 -7328
rect 8372 -7582 8468 -7486
<< metal2 >>
rect 5042 1080 5138 1090
rect 5042 974 5138 984
rect 5876 824 5946 834
rect 5876 700 5946 764
rect 7504 820 7564 830
rect 5870 694 5946 700
rect 5996 694 6036 754
rect 6096 694 6166 754
rect 6226 694 6316 754
rect 6376 694 6446 754
rect 6506 694 6566 754
rect 6886 694 6926 754
rect 6986 694 7056 754
rect 7116 694 7206 754
rect 7266 694 7336 754
rect 7396 694 7456 754
rect 7504 710 7564 760
rect 7503 700 7572 710
rect 5870 684 5876 694
rect 5866 634 5876 684
rect 5866 624 5946 634
rect 5870 458 5930 624
rect 6166 602 6226 694
rect 7040 604 7100 694
rect 7503 621 7572 631
rect 6159 546 6168 602
rect 6224 546 6233 602
rect 7033 548 7042 604
rect 7098 548 7107 604
rect 7040 546 7100 548
rect 6166 544 6226 546
rect 5863 402 5872 458
rect 5928 402 5937 458
rect 5870 400 5930 402
rect 7504 372 7564 621
rect 8416 536 8512 546
rect 8416 430 8512 440
rect 7504 316 7506 372
rect 7562 316 7564 372
rect 7504 314 7564 316
rect 7506 307 7562 314
rect 6130 208 7170 210
rect 6123 152 6132 208
rect 6188 152 7170 208
rect 6130 150 7170 152
rect 7230 150 7239 210
rect 6000 118 7040 120
rect 5993 62 6002 118
rect 6058 62 7040 118
rect 6000 60 7040 62
rect 7100 60 7109 120
rect 5870 28 6910 30
rect 5863 -28 5872 28
rect 5928 -28 6910 28
rect 5870 -30 6910 -28
rect 6970 -30 6979 30
rect 5740 -62 6780 -60
rect 5733 -118 5742 -62
rect 5798 -118 6780 -62
rect 5740 -120 6780 -118
rect 6840 -120 6849 -60
rect 5062 -160 5158 -150
rect 5062 -266 5158 -256
rect 6392 -482 6448 -475
rect 6034 -484 6190 -482
rect 6308 -484 6450 -482
rect 6780 -484 6910 -482
rect 5863 -546 5872 -490
rect 5928 -546 5937 -490
rect 6034 -540 6132 -484
rect 6188 -540 6197 -484
rect 6308 -540 6392 -484
rect 6448 -540 6450 -484
rect 6034 -542 6190 -540
rect 6308 -542 6450 -540
rect 6643 -542 6652 -486
rect 6708 -542 6717 -486
rect 6773 -540 6782 -484
rect 6838 -540 6910 -484
rect 6780 -542 6910 -540
rect 6392 -549 6448 -542
rect 7033 -552 7042 -496
rect 7098 -552 7107 -496
rect 7293 -546 7302 -490
rect 7358 -546 7367 -490
rect 7620 -564 7680 -482
rect 7560 -566 7680 -564
rect 7553 -622 7562 -566
rect 7618 -622 7680 -566
rect 7560 -624 7680 -622
rect 8386 -704 8482 -694
rect 8386 -810 8482 -800
rect 5032 -960 5128 -950
rect 5032 -1066 5128 -1056
rect 6306 -1288 6450 -1286
rect 6652 -1288 6708 -1279
rect 6038 -1290 6190 -1288
rect 5740 -1292 5912 -1290
rect 5733 -1348 5742 -1292
rect 5798 -1348 5912 -1292
rect 6038 -1346 6132 -1290
rect 6188 -1346 6197 -1290
rect 6306 -1344 6392 -1288
rect 6448 -1344 6457 -1288
rect 6306 -1346 6450 -1344
rect 6038 -1348 6190 -1346
rect 5740 -1350 5912 -1348
rect 6652 -1353 6708 -1344
rect 6848 -1292 6970 -1290
rect 6848 -1348 6912 -1292
rect 6968 -1348 6977 -1292
rect 7033 -1342 7042 -1286
rect 7098 -1342 7107 -1286
rect 7293 -1346 7302 -1290
rect 7358 -1346 7367 -1290
rect 6848 -1350 6970 -1348
rect 7614 -1382 7674 -1290
rect 7560 -1384 7674 -1382
rect 7553 -1440 7562 -1384
rect 7618 -1440 7674 -1384
rect 7560 -1442 7674 -1440
rect 8398 -1504 8494 -1494
rect 8398 -1610 8494 -1600
rect 5052 -1760 5148 -1750
rect 5052 -1866 5148 -1856
rect 5863 -2142 5872 -2086
rect 5928 -2142 5937 -2086
rect 6324 -2088 6450 -2086
rect 5993 -2148 6002 -2092
rect 6058 -2148 6067 -2092
rect 6324 -2144 6392 -2088
rect 6448 -2144 6457 -2088
rect 6643 -2138 6652 -2082
rect 6708 -2138 6717 -2082
rect 6780 -2092 6906 -2090
rect 6324 -2146 6450 -2144
rect 6773 -2148 6782 -2092
rect 6838 -2148 6906 -2092
rect 6780 -2150 6906 -2148
rect 7032 -2094 7230 -2092
rect 7032 -2150 7172 -2094
rect 7228 -2150 7237 -2094
rect 7293 -2144 7302 -2088
rect 7358 -2144 7367 -2088
rect 7032 -2152 7230 -2150
rect 7614 -2166 7674 -2100
rect 7560 -2168 7674 -2166
rect 7553 -2224 7562 -2168
rect 7618 -2224 7674 -2168
rect 7560 -2226 7674 -2224
rect 8396 -2304 8492 -2294
rect 8396 -2410 8492 -2400
rect 5046 -2559 5142 -2549
rect 5046 -2665 5142 -2655
rect 5740 -2884 5904 -2882
rect 5733 -2940 5742 -2884
rect 5798 -2940 5904 -2884
rect 5740 -2942 5904 -2940
rect 5993 -2942 6002 -2886
rect 6058 -2942 6067 -2886
rect 6320 -2890 6450 -2888
rect 6320 -2946 6392 -2890
rect 6448 -2946 6457 -2890
rect 6643 -2944 6652 -2888
rect 6708 -2944 6717 -2888
rect 6850 -2892 6970 -2890
rect 6320 -2948 6450 -2946
rect 6850 -2948 6912 -2892
rect 6968 -2948 6977 -2892
rect 7026 -2898 7230 -2896
rect 6850 -2950 6970 -2948
rect 7026 -2954 7172 -2898
rect 7228 -2954 7237 -2898
rect 7293 -2940 7302 -2884
rect 7358 -2940 7367 -2884
rect 7026 -2956 7230 -2954
rect 7620 -2980 7680 -2888
rect 7560 -2982 7680 -2980
rect 7553 -3038 7562 -2982
rect 7618 -3038 7680 -2982
rect 7560 -3040 7680 -3038
rect 8380 -3104 8476 -3094
rect 8380 -3210 8476 -3200
rect 5062 -3360 5158 -3350
rect 5062 -3466 5158 -3456
rect 5863 -3740 5872 -3684
rect 5928 -3740 5937 -3684
rect 6054 -3688 6190 -3686
rect 6054 -3744 6132 -3688
rect 6188 -3744 6197 -3688
rect 6253 -3740 6262 -3684
rect 6318 -3740 6327 -3684
rect 6054 -3746 6190 -3744
rect 6643 -3746 6652 -3690
rect 6708 -3746 6717 -3690
rect 6780 -3694 6906 -3692
rect 6773 -3750 6782 -3694
rect 6838 -3750 6906 -3694
rect 6780 -3752 6906 -3750
rect 7033 -3754 7042 -3698
rect 7098 -3754 7107 -3698
rect 7304 -3770 7364 -3694
rect 7432 -3770 7488 -3763
rect 7304 -3772 7490 -3770
rect 7304 -3828 7432 -3772
rect 7488 -3828 7490 -3772
rect 7618 -3774 7678 -3682
rect 7560 -3776 7678 -3774
rect 7304 -3830 7490 -3828
rect 7432 -3837 7488 -3830
rect 7553 -3832 7562 -3776
rect 7618 -3832 7678 -3776
rect 7560 -3834 7678 -3832
rect 8370 -3904 8466 -3894
rect 8370 -4010 8466 -4000
rect 5036 -4160 5132 -4150
rect 5036 -4266 5132 -4256
rect 6052 -4488 6190 -4486
rect 5740 -4496 5916 -4494
rect 5733 -4552 5742 -4496
rect 5798 -4552 5916 -4496
rect 6052 -4544 6132 -4488
rect 6188 -4544 6197 -4488
rect 6052 -4546 6190 -4544
rect 6253 -4548 6262 -4492
rect 6318 -4548 6327 -4492
rect 6643 -4542 6652 -4486
rect 6708 -4542 6717 -4486
rect 6858 -4488 6970 -4486
rect 6858 -4544 6912 -4488
rect 6968 -4544 6977 -4488
rect 7033 -4542 7042 -4486
rect 7098 -4542 7107 -4486
rect 6858 -4546 6970 -4544
rect 5740 -4554 5916 -4552
rect 7298 -4572 7358 -4492
rect 7432 -4572 7488 -4565
rect 7616 -4570 7676 -4486
rect 7560 -4572 7676 -4570
rect 7298 -4574 7490 -4572
rect 7298 -4630 7432 -4574
rect 7488 -4630 7490 -4574
rect 7553 -4628 7562 -4572
rect 7618 -4628 7676 -4572
rect 7560 -4630 7676 -4628
rect 7298 -4632 7490 -4630
rect 7432 -4639 7488 -4632
rect 8388 -4704 8484 -4694
rect 8388 -4810 8484 -4800
rect 5036 -4960 5132 -4950
rect 5036 -5066 5132 -5056
rect 5863 -5346 5872 -5290
rect 5928 -5346 5937 -5290
rect 6780 -5292 6902 -5290
rect 5993 -5348 6002 -5292
rect 6058 -5348 6067 -5292
rect 6253 -5350 6262 -5294
rect 6318 -5350 6327 -5294
rect 6643 -5348 6652 -5292
rect 6708 -5348 6717 -5292
rect 6773 -5348 6782 -5292
rect 6838 -5348 6902 -5292
rect 6780 -5350 6902 -5348
rect 7032 -5296 7230 -5294
rect 7032 -5352 7172 -5296
rect 7228 -5352 7237 -5296
rect 7032 -5354 7230 -5352
rect 7314 -5382 7374 -5296
rect 7620 -5380 7680 -5288
rect 7560 -5382 7680 -5380
rect 7314 -5384 7490 -5382
rect 7314 -5440 7432 -5384
rect 7488 -5440 7497 -5384
rect 7553 -5438 7562 -5382
rect 7618 -5438 7680 -5382
rect 7560 -5440 7680 -5438
rect 7314 -5442 7490 -5440
rect 8370 -5504 8466 -5494
rect 8370 -5610 8466 -5600
rect 5032 -5760 5128 -5750
rect 5032 -5866 5128 -5856
rect 7022 -6082 7230 -6080
rect 5740 -6102 5908 -6100
rect 5733 -6158 5742 -6102
rect 5798 -6158 5908 -6102
rect 5993 -6146 6002 -6090
rect 6058 -6146 6067 -6090
rect 6253 -6146 6262 -6090
rect 6318 -6146 6327 -6090
rect 6643 -6142 6652 -6086
rect 6708 -6142 6717 -6086
rect 6838 -6090 6970 -6088
rect 6838 -6146 6912 -6090
rect 6968 -6146 6977 -6090
rect 7022 -6138 7172 -6082
rect 7228 -6138 7237 -6082
rect 7022 -6140 7230 -6138
rect 6838 -6148 6970 -6146
rect 5740 -6160 5908 -6158
rect 7304 -6176 7364 -6090
rect 7304 -6178 7490 -6176
rect 7304 -6234 7432 -6178
rect 7488 -6234 7497 -6178
rect 7618 -6180 7678 -6094
rect 7560 -6182 7678 -6180
rect 7304 -6236 7490 -6234
rect 7553 -6238 7562 -6182
rect 7618 -6238 7678 -6182
rect 7560 -6240 7678 -6238
rect 8394 -6303 8490 -6293
rect 8394 -6409 8490 -6399
rect 6260 -6452 7300 -6450
rect 6253 -6508 6262 -6452
rect 6318 -6508 7300 -6452
rect 6260 -6510 7300 -6508
rect 7360 -6510 7369 -6450
rect 6390 -6542 7430 -6540
rect 6383 -6598 6392 -6542
rect 6448 -6598 7430 -6542
rect 6390 -6600 7430 -6598
rect 7490 -6600 7499 -6540
rect 6520 -6632 7560 -6630
rect 6513 -6688 6522 -6632
rect 6578 -6688 7560 -6632
rect 6520 -6690 7560 -6688
rect 7620 -6690 7629 -6630
rect 6650 -6722 7690 -6720
rect 6643 -6778 6652 -6722
rect 6708 -6778 7690 -6722
rect 6650 -6780 7690 -6778
rect 7750 -6780 7759 -6720
rect 5032 -6948 5128 -6938
rect 7158 -7002 7214 -6995
rect 5032 -7054 5128 -7044
rect 7156 -7004 7216 -7002
rect 6634 -7052 6694 -7050
rect 6260 -7058 6320 -7056
rect 6253 -7114 6262 -7058
rect 6318 -7114 6327 -7058
rect 6627 -7108 6636 -7052
rect 6692 -7108 6701 -7052
rect 7156 -7060 7158 -7004
rect 7214 -7060 7216 -7004
rect 6260 -7260 6320 -7114
rect 6634 -7200 6694 -7108
rect 6025 -7320 6065 -7260
rect 6125 -7320 6195 -7260
rect 6255 -7320 6345 -7260
rect 6405 -7320 6475 -7260
rect 6535 -7320 6595 -7260
rect 6634 -7328 6694 -7260
rect 7156 -7264 7216 -7060
rect 7534 -7198 7594 -7194
rect 7534 -7200 7750 -7198
rect 7594 -7256 7692 -7200
rect 7748 -7256 7757 -7200
rect 7594 -7258 7750 -7256
rect 6913 -7324 6953 -7264
rect 7013 -7324 7083 -7264
rect 7143 -7324 7233 -7264
rect 7293 -7324 7363 -7264
rect 7423 -7324 7483 -7264
rect 6634 -7394 6694 -7388
rect 7534 -7328 7594 -7260
rect 7534 -7394 7594 -7388
rect 8372 -7486 8468 -7476
rect 8372 -7592 8468 -7582
<< via2 >>
rect 5042 984 5138 1080
rect 6168 546 6224 602
rect 7042 548 7098 604
rect 5872 402 5928 458
rect 8416 440 8512 536
rect 7506 316 7562 372
rect 6132 152 6188 208
rect 7170 150 7230 210
rect 6002 62 6058 118
rect 7040 60 7100 120
rect 5872 -28 5928 28
rect 6910 -30 6970 30
rect 5742 -118 5798 -62
rect 6780 -120 6840 -60
rect 5062 -256 5158 -160
rect 5872 -546 5928 -490
rect 6132 -540 6188 -484
rect 6392 -540 6448 -484
rect 6652 -542 6708 -486
rect 6782 -540 6838 -484
rect 7042 -552 7098 -496
rect 7302 -546 7358 -490
rect 7562 -622 7618 -566
rect 8386 -800 8482 -704
rect 5032 -1056 5128 -960
rect 5742 -1348 5798 -1292
rect 6132 -1346 6188 -1290
rect 6392 -1344 6448 -1288
rect 6652 -1344 6708 -1288
rect 6912 -1348 6968 -1292
rect 7042 -1342 7098 -1286
rect 7302 -1346 7358 -1290
rect 7562 -1440 7618 -1384
rect 8398 -1600 8494 -1504
rect 5052 -1856 5148 -1760
rect 5872 -2142 5928 -2086
rect 6002 -2148 6058 -2092
rect 6392 -2144 6448 -2088
rect 6652 -2138 6708 -2082
rect 6782 -2148 6838 -2092
rect 7172 -2150 7228 -2094
rect 7302 -2144 7358 -2088
rect 7562 -2224 7618 -2168
rect 8396 -2400 8492 -2304
rect 5046 -2655 5142 -2559
rect 5742 -2940 5798 -2884
rect 6002 -2942 6058 -2886
rect 6392 -2946 6448 -2890
rect 6652 -2944 6708 -2888
rect 6912 -2948 6968 -2892
rect 7172 -2954 7228 -2898
rect 7302 -2940 7358 -2884
rect 7562 -3038 7618 -2982
rect 8380 -3200 8476 -3104
rect 5062 -3456 5158 -3360
rect 5872 -3740 5928 -3684
rect 6132 -3744 6188 -3688
rect 6262 -3740 6318 -3684
rect 6652 -3746 6708 -3690
rect 6782 -3750 6838 -3694
rect 7042 -3754 7098 -3698
rect 7432 -3828 7488 -3772
rect 7562 -3832 7618 -3776
rect 8370 -4000 8466 -3904
rect 5036 -4256 5132 -4160
rect 5742 -4552 5798 -4496
rect 6132 -4544 6188 -4488
rect 6262 -4548 6318 -4492
rect 6652 -4542 6708 -4486
rect 6912 -4544 6968 -4488
rect 7042 -4542 7098 -4486
rect 7432 -4630 7488 -4574
rect 7562 -4628 7618 -4572
rect 8388 -4800 8484 -4704
rect 5036 -5056 5132 -4960
rect 5872 -5346 5928 -5290
rect 6002 -5348 6058 -5292
rect 6262 -5350 6318 -5294
rect 6652 -5348 6708 -5292
rect 6782 -5348 6838 -5292
rect 7172 -5352 7228 -5296
rect 7432 -5440 7488 -5384
rect 7562 -5438 7618 -5382
rect 8370 -5600 8466 -5504
rect 5032 -5856 5128 -5760
rect 5742 -6158 5798 -6102
rect 6002 -6146 6058 -6090
rect 6262 -6146 6318 -6090
rect 6652 -6142 6708 -6086
rect 6912 -6146 6968 -6090
rect 7172 -6138 7228 -6082
rect 7432 -6234 7488 -6178
rect 7562 -6238 7618 -6182
rect 8394 -6399 8490 -6303
rect 6262 -6508 6318 -6452
rect 7300 -6510 7360 -6450
rect 6392 -6598 6448 -6542
rect 7430 -6600 7490 -6540
rect 6522 -6688 6578 -6632
rect 7560 -6690 7620 -6630
rect 6652 -6778 6708 -6722
rect 7690 -6780 7750 -6720
rect 5032 -7044 5128 -6948
rect 6262 -7114 6318 -7058
rect 6636 -7108 6692 -7052
rect 7158 -7060 7214 -7004
rect 7692 -7256 7748 -7200
rect 8372 -7582 8468 -7486
<< metal3 >>
rect 5032 1080 5148 1085
rect 5032 984 5042 1080
rect 5138 984 5148 1080
rect 5032 979 5148 984
rect 6163 604 6229 607
rect 5740 602 6229 604
rect 5740 546 6168 602
rect 6224 546 6229 602
rect 5740 544 6229 546
rect 5740 -57 5800 544
rect 6163 541 6229 544
rect 7037 604 7103 609
rect 7037 548 7042 604
rect 7098 548 7103 604
rect 7037 543 7103 548
rect 5867 458 5933 463
rect 5867 402 5872 458
rect 5928 402 5933 458
rect 5867 397 5933 402
rect 5870 33 5930 397
rect 6000 123 6060 324
rect 6130 213 6190 324
rect 6127 208 6193 213
rect 6127 152 6132 208
rect 6188 152 6193 208
rect 6127 147 6193 152
rect 5997 118 6063 123
rect 5997 62 6002 118
rect 6058 62 6063 118
rect 5997 57 6063 62
rect 5867 28 5933 33
rect 5867 -28 5872 28
rect 5928 -28 5933 28
rect 5867 -33 5933 -28
rect 5737 -62 5803 -57
rect 5737 -118 5742 -62
rect 5798 -118 5803 -62
rect 5737 -123 5803 -118
rect 5052 -160 5168 -155
rect 5052 -256 5062 -160
rect 5158 -256 5168 -160
rect 5052 -261 5168 -256
rect 5022 -960 5138 -955
rect 5022 -1056 5032 -960
rect 5128 -1056 5138 -960
rect 5022 -1061 5138 -1056
rect 5740 -1287 5800 -123
rect 5870 -485 5930 -33
rect 5867 -490 5933 -485
rect 5867 -546 5872 -490
rect 5928 -546 5933 -490
rect 5867 -551 5933 -546
rect 5737 -1292 5803 -1287
rect 5737 -1348 5742 -1292
rect 5798 -1348 5803 -1292
rect 5737 -1353 5803 -1348
rect 5042 -1760 5158 -1755
rect 5042 -1856 5052 -1760
rect 5148 -1856 5158 -1760
rect 5042 -1861 5158 -1856
rect 5036 -2559 5152 -2554
rect 5036 -2655 5046 -2559
rect 5142 -2655 5152 -2559
rect 5036 -2660 5152 -2655
rect 5740 -2879 5800 -1353
rect 5870 -2081 5930 -551
rect 5867 -2086 5933 -2081
rect 5867 -2142 5872 -2086
rect 5928 -2142 5933 -2086
rect 6000 -2087 6060 57
rect 6130 -479 6190 147
rect 6127 -484 6193 -479
rect 6127 -540 6132 -484
rect 6188 -540 6193 -484
rect 6127 -545 6193 -540
rect 6130 -1285 6190 -545
rect 6127 -1290 6193 -1285
rect 6127 -1346 6132 -1290
rect 6188 -1346 6193 -1290
rect 6127 -1351 6193 -1346
rect 5867 -2147 5933 -2142
rect 5997 -2092 6063 -2087
rect 5737 -2884 5803 -2879
rect 5737 -2940 5742 -2884
rect 5798 -2940 5803 -2884
rect 5737 -2945 5803 -2940
rect 5052 -3360 5168 -3355
rect 5052 -3456 5062 -3360
rect 5158 -3456 5168 -3360
rect 5052 -3461 5168 -3456
rect 5026 -4160 5142 -4155
rect 5026 -4256 5036 -4160
rect 5132 -4256 5142 -4160
rect 5026 -4261 5142 -4256
rect 5740 -4491 5800 -2945
rect 5870 -3679 5930 -2147
rect 5997 -2148 6002 -2092
rect 6058 -2148 6063 -2092
rect 5997 -2153 6063 -2148
rect 6000 -2881 6060 -2153
rect 5997 -2886 6063 -2881
rect 5997 -2942 6002 -2886
rect 6058 -2942 6063 -2886
rect 5997 -2947 6063 -2942
rect 5867 -3684 5933 -3679
rect 5867 -3740 5872 -3684
rect 5928 -3740 5933 -3684
rect 5867 -3745 5933 -3740
rect 5737 -4496 5803 -4491
rect 5737 -4552 5742 -4496
rect 5798 -4552 5803 -4496
rect 5737 -4557 5803 -4552
rect 5026 -4960 5142 -4955
rect 5026 -5056 5036 -4960
rect 5132 -5056 5142 -4960
rect 5026 -5061 5142 -5056
rect 5022 -5760 5138 -5755
rect 5022 -5856 5032 -5760
rect 5128 -5856 5138 -5760
rect 5022 -5861 5138 -5856
rect 5740 -6097 5800 -4557
rect 5870 -5285 5930 -3745
rect 5867 -5290 5933 -5285
rect 6000 -5287 6060 -2947
rect 6130 -3683 6190 -1351
rect 6260 -3679 6320 324
rect 6390 -479 6450 324
rect 6387 -484 6453 -479
rect 6387 -540 6392 -484
rect 6448 -540 6453 -484
rect 6387 -545 6453 -540
rect 6390 -1283 6450 -545
rect 6387 -1288 6453 -1283
rect 6387 -1344 6392 -1288
rect 6448 -1344 6453 -1288
rect 6387 -1349 6453 -1344
rect 6390 -2083 6450 -1349
rect 6387 -2088 6453 -2083
rect 6387 -2144 6392 -2088
rect 6448 -2144 6453 -2088
rect 6387 -2149 6453 -2144
rect 6390 -2885 6450 -2149
rect 6387 -2890 6453 -2885
rect 6387 -2946 6392 -2890
rect 6448 -2946 6453 -2890
rect 6387 -2951 6453 -2946
rect 6127 -3688 6193 -3683
rect 6127 -3744 6132 -3688
rect 6188 -3744 6193 -3688
rect 6127 -3749 6193 -3744
rect 6257 -3684 6323 -3679
rect 6257 -3740 6262 -3684
rect 6318 -3740 6323 -3684
rect 6257 -3745 6323 -3740
rect 6130 -4483 6190 -3749
rect 6127 -4488 6193 -4483
rect 6260 -4487 6320 -3745
rect 6127 -4544 6132 -4488
rect 6188 -4544 6193 -4488
rect 6127 -4549 6193 -4544
rect 6257 -4492 6323 -4487
rect 6257 -4548 6262 -4492
rect 6318 -4548 6323 -4492
rect 5867 -5346 5872 -5290
rect 5928 -5346 5933 -5290
rect 5867 -5351 5933 -5346
rect 5997 -5292 6063 -5287
rect 5997 -5348 6002 -5292
rect 6058 -5348 6063 -5292
rect 5737 -6102 5803 -6097
rect 5737 -6158 5742 -6102
rect 5798 -6158 5803 -6102
rect 5737 -6163 5803 -6158
rect 5740 -6460 5800 -6163
rect 5870 -6460 5930 -5351
rect 5997 -5353 6063 -5348
rect 6000 -6085 6060 -5353
rect 5997 -6090 6063 -6085
rect 5997 -6146 6002 -6090
rect 6058 -6146 6063 -6090
rect 5997 -6151 6063 -6146
rect 6000 -6460 6060 -6151
rect 6130 -6460 6190 -4549
rect 6257 -4553 6323 -4548
rect 6260 -5289 6320 -4553
rect 6257 -5294 6323 -5289
rect 6257 -5350 6262 -5294
rect 6318 -5350 6323 -5294
rect 6257 -5355 6323 -5350
rect 6260 -6085 6320 -5355
rect 6257 -6090 6323 -6085
rect 6257 -6146 6262 -6090
rect 6318 -6146 6323 -6090
rect 6257 -6151 6323 -6146
rect 6260 -6447 6320 -6151
rect 6257 -6452 6323 -6447
rect 6257 -6508 6262 -6452
rect 6318 -6508 6323 -6452
rect 6257 -6513 6323 -6508
rect 5022 -6948 5138 -6943
rect 5022 -7044 5032 -6948
rect 5128 -7044 5138 -6948
rect 5022 -7049 5138 -7044
rect 6260 -7053 6320 -6513
rect 6390 -6537 6450 -2951
rect 6387 -6542 6453 -6537
rect 6387 -6598 6392 -6542
rect 6448 -6598 6453 -6542
rect 6387 -6603 6453 -6598
rect 6390 -7050 6450 -6603
rect 6520 -6627 6580 324
rect 6650 -481 6710 324
rect 6780 -55 6840 250
rect 6910 35 6970 250
rect 7040 125 7100 543
rect 8406 536 8522 541
rect 8406 440 8416 536
rect 8512 440 8522 536
rect 8406 435 8522 440
rect 7501 374 7567 377
rect 7170 372 7567 374
rect 7170 316 7506 372
rect 7562 316 7567 372
rect 7170 314 7567 316
rect 7170 215 7230 314
rect 7501 311 7567 314
rect 7165 210 7235 215
rect 7165 150 7170 210
rect 7230 150 7235 210
rect 7165 145 7235 150
rect 7035 120 7105 125
rect 7035 60 7040 120
rect 7100 60 7105 120
rect 7035 55 7105 60
rect 6905 30 6975 35
rect 6905 -30 6910 30
rect 6970 -30 6975 30
rect 6905 -35 6975 -30
rect 6775 -60 6845 -55
rect 6775 -120 6780 -60
rect 6840 -120 6845 -60
rect 6775 -125 6845 -120
rect 6780 -479 6840 -125
rect 6647 -486 6713 -481
rect 6647 -542 6652 -486
rect 6708 -542 6713 -486
rect 6647 -547 6713 -542
rect 6777 -484 6843 -479
rect 6777 -540 6782 -484
rect 6838 -540 6843 -484
rect 6777 -545 6843 -540
rect 6650 -1283 6710 -547
rect 6647 -1288 6713 -1283
rect 6647 -1344 6652 -1288
rect 6708 -1344 6713 -1288
rect 6647 -1349 6713 -1344
rect 6650 -2077 6710 -1349
rect 6647 -2082 6713 -2077
rect 6647 -2138 6652 -2082
rect 6708 -2138 6713 -2082
rect 6780 -2087 6840 -545
rect 6910 -1287 6970 -35
rect 7040 -491 7100 55
rect 7037 -496 7103 -491
rect 7037 -552 7042 -496
rect 7098 -552 7103 -496
rect 7037 -557 7103 -552
rect 7040 -1281 7100 -557
rect 7037 -1286 7103 -1281
rect 6907 -1292 6973 -1287
rect 6907 -1348 6912 -1292
rect 6968 -1348 6973 -1292
rect 7037 -1342 7042 -1286
rect 7098 -1342 7103 -1286
rect 7037 -1347 7103 -1342
rect 6907 -1353 6973 -1348
rect 6647 -2143 6713 -2138
rect 6777 -2092 6843 -2087
rect 6650 -2883 6710 -2143
rect 6777 -2148 6782 -2092
rect 6838 -2148 6843 -2092
rect 6777 -2153 6843 -2148
rect 6647 -2888 6713 -2883
rect 6647 -2944 6652 -2888
rect 6708 -2944 6713 -2888
rect 6647 -2949 6713 -2944
rect 6650 -3685 6710 -2949
rect 6647 -3690 6713 -3685
rect 6780 -3689 6840 -2153
rect 6910 -2887 6970 -1353
rect 6907 -2892 6973 -2887
rect 6907 -2948 6912 -2892
rect 6968 -2948 6973 -2892
rect 6907 -2953 6973 -2948
rect 6647 -3746 6652 -3690
rect 6708 -3746 6713 -3690
rect 6647 -3751 6713 -3746
rect 6777 -3694 6843 -3689
rect 6777 -3750 6782 -3694
rect 6838 -3750 6843 -3694
rect 6650 -4481 6710 -3751
rect 6777 -3755 6843 -3750
rect 6647 -4486 6713 -4481
rect 6647 -4542 6652 -4486
rect 6708 -4542 6713 -4486
rect 6647 -4547 6713 -4542
rect 6650 -5287 6710 -4547
rect 6780 -5287 6840 -3755
rect 6910 -4483 6970 -2953
rect 7040 -3693 7100 -1347
rect 7170 -2089 7230 145
rect 7300 -485 7360 -90
rect 7297 -490 7363 -485
rect 7297 -546 7302 -490
rect 7358 -546 7363 -490
rect 7297 -551 7363 -546
rect 7300 -1285 7360 -551
rect 7297 -1290 7363 -1285
rect 7297 -1346 7302 -1290
rect 7358 -1346 7363 -1290
rect 7297 -1351 7363 -1346
rect 7300 -2083 7360 -1351
rect 7297 -2088 7363 -2083
rect 7167 -2094 7233 -2089
rect 7167 -2150 7172 -2094
rect 7228 -2150 7233 -2094
rect 7297 -2144 7302 -2088
rect 7358 -2144 7363 -2088
rect 7297 -2149 7363 -2144
rect 7167 -2155 7233 -2150
rect 7170 -2893 7230 -2155
rect 7300 -2879 7360 -2149
rect 7297 -2884 7363 -2879
rect 7167 -2898 7233 -2893
rect 7167 -2954 7172 -2898
rect 7228 -2954 7233 -2898
rect 7297 -2940 7302 -2884
rect 7358 -2940 7363 -2884
rect 7297 -2945 7363 -2940
rect 7167 -2959 7233 -2954
rect 7037 -3698 7103 -3693
rect 7037 -3754 7042 -3698
rect 7098 -3754 7103 -3698
rect 7037 -3759 7103 -3754
rect 7040 -4481 7100 -3759
rect 6907 -4488 6973 -4483
rect 6907 -4544 6912 -4488
rect 6968 -4544 6973 -4488
rect 6907 -4549 6973 -4544
rect 7037 -4486 7103 -4481
rect 7037 -4542 7042 -4486
rect 7098 -4542 7103 -4486
rect 7037 -4547 7103 -4542
rect 6647 -5292 6713 -5287
rect 6647 -5348 6652 -5292
rect 6708 -5348 6713 -5292
rect 6647 -5353 6713 -5348
rect 6777 -5292 6843 -5287
rect 6777 -5348 6782 -5292
rect 6838 -5348 6843 -5292
rect 6777 -5353 6843 -5348
rect 6650 -6081 6710 -5353
rect 6647 -6086 6713 -6081
rect 6647 -6142 6652 -6086
rect 6708 -6142 6713 -6086
rect 6647 -6147 6713 -6142
rect 6517 -6632 6583 -6627
rect 6517 -6688 6522 -6632
rect 6578 -6688 6583 -6632
rect 6517 -6693 6583 -6688
rect 6520 -6830 6580 -6693
rect 6650 -6717 6710 -6147
rect 6647 -6722 6713 -6717
rect 6647 -6778 6652 -6722
rect 6708 -6778 6713 -6722
rect 6647 -6783 6713 -6778
rect 6650 -6830 6710 -6783
rect 6780 -6830 6840 -5353
rect 6910 -6085 6970 -4549
rect 6907 -6090 6973 -6085
rect 6907 -6146 6912 -6090
rect 6968 -6146 6973 -6090
rect 6907 -6151 6973 -6146
rect 6910 -6830 6970 -6151
rect 7040 -6830 7100 -4547
rect 7170 -5291 7230 -2959
rect 7167 -5296 7233 -5291
rect 7167 -5352 7172 -5296
rect 7228 -5352 7233 -5296
rect 7167 -5357 7233 -5352
rect 7170 -6077 7230 -5357
rect 7167 -6082 7233 -6077
rect 7167 -6138 7172 -6082
rect 7228 -6138 7233 -6082
rect 7167 -6143 7233 -6138
rect 7170 -6830 7230 -6143
rect 7300 -6445 7360 -2945
rect 7430 -3767 7490 -90
rect 7560 -561 7620 -90
rect 7557 -566 7623 -561
rect 7557 -622 7562 -566
rect 7618 -622 7623 -566
rect 7557 -627 7623 -622
rect 7560 -1379 7620 -627
rect 7557 -1384 7623 -1379
rect 7557 -1440 7562 -1384
rect 7618 -1440 7623 -1384
rect 7557 -1445 7623 -1440
rect 7560 -2163 7620 -1445
rect 7557 -2168 7623 -2163
rect 7557 -2224 7562 -2168
rect 7618 -2224 7623 -2168
rect 7557 -2229 7623 -2224
rect 7560 -2977 7620 -2229
rect 7557 -2982 7623 -2977
rect 7557 -3038 7562 -2982
rect 7618 -3038 7623 -2982
rect 7557 -3043 7623 -3038
rect 7427 -3772 7493 -3767
rect 7560 -3771 7620 -3043
rect 7427 -3828 7432 -3772
rect 7488 -3828 7493 -3772
rect 7427 -3833 7493 -3828
rect 7557 -3776 7623 -3771
rect 7557 -3832 7562 -3776
rect 7618 -3832 7623 -3776
rect 7430 -4569 7490 -3833
rect 7557 -3837 7623 -3832
rect 7560 -4567 7620 -3837
rect 7427 -4574 7493 -4569
rect 7427 -4630 7432 -4574
rect 7488 -4630 7493 -4574
rect 7427 -4635 7493 -4630
rect 7557 -4572 7623 -4567
rect 7557 -4628 7562 -4572
rect 7618 -4628 7623 -4572
rect 7557 -4633 7623 -4628
rect 7430 -5379 7490 -4635
rect 7560 -5377 7620 -4633
rect 7427 -5384 7493 -5379
rect 7427 -5440 7432 -5384
rect 7488 -5440 7493 -5384
rect 7427 -5445 7493 -5440
rect 7557 -5382 7623 -5377
rect 7557 -5438 7562 -5382
rect 7618 -5438 7623 -5382
rect 7557 -5443 7623 -5438
rect 7430 -6173 7490 -5445
rect 7427 -6178 7493 -6173
rect 7560 -6177 7620 -5443
rect 7427 -6234 7432 -6178
rect 7488 -6234 7493 -6178
rect 7427 -6239 7493 -6234
rect 7557 -6182 7623 -6177
rect 7557 -6238 7562 -6182
rect 7618 -6238 7623 -6182
rect 7295 -6450 7365 -6445
rect 7295 -6510 7300 -6450
rect 7360 -6510 7365 -6450
rect 7295 -6515 7365 -6510
rect 7300 -6830 7360 -6515
rect 7430 -6535 7490 -6239
rect 7557 -6243 7623 -6238
rect 7425 -6540 7495 -6535
rect 7425 -6600 7430 -6540
rect 7490 -6600 7495 -6540
rect 7425 -6605 7495 -6600
rect 7430 -6830 7490 -6605
rect 7560 -6625 7620 -6243
rect 7555 -6630 7625 -6625
rect 7555 -6690 7560 -6630
rect 7620 -6690 7625 -6630
rect 7555 -6695 7625 -6690
rect 7153 -7002 7219 -6999
rect 7560 -7002 7620 -6695
rect 7690 -6715 7750 -90
rect 8376 -704 8492 -699
rect 8376 -800 8386 -704
rect 8482 -800 8492 -704
rect 8376 -805 8492 -800
rect 8388 -1504 8504 -1499
rect 8388 -1600 8398 -1504
rect 8494 -1600 8504 -1504
rect 8388 -1605 8504 -1600
rect 8386 -2304 8502 -2299
rect 8386 -2400 8396 -2304
rect 8492 -2400 8502 -2304
rect 8386 -2405 8502 -2400
rect 8370 -3104 8486 -3099
rect 8370 -3200 8380 -3104
rect 8476 -3200 8486 -3104
rect 8370 -3205 8486 -3200
rect 8360 -3904 8476 -3899
rect 8360 -4000 8370 -3904
rect 8466 -4000 8476 -3904
rect 8360 -4005 8476 -4000
rect 8378 -4704 8494 -4699
rect 8378 -4800 8388 -4704
rect 8484 -4800 8494 -4704
rect 8378 -4805 8494 -4800
rect 8360 -5504 8476 -5499
rect 8360 -5600 8370 -5504
rect 8466 -5600 8476 -5504
rect 8360 -5605 8476 -5600
rect 8384 -6303 8500 -6298
rect 8384 -6399 8394 -6303
rect 8490 -6399 8500 -6303
rect 8384 -6404 8500 -6399
rect 7685 -6720 7755 -6715
rect 7685 -6780 7690 -6720
rect 7750 -6780 7755 -6720
rect 7685 -6785 7755 -6780
rect 7153 -7004 7620 -7002
rect 6631 -7050 6697 -7047
rect 6390 -7052 6697 -7050
rect 6257 -7058 6323 -7053
rect 6257 -7114 6262 -7058
rect 6318 -7114 6323 -7058
rect 6390 -7108 6636 -7052
rect 6692 -7108 6697 -7052
rect 7153 -7060 7158 -7004
rect 7214 -7060 7620 -7004
rect 7153 -7062 7620 -7060
rect 7153 -7065 7219 -7062
rect 6390 -7110 6697 -7108
rect 6631 -7113 6697 -7110
rect 6257 -7119 6323 -7114
rect 7690 -7195 7750 -6785
rect 7687 -7200 7753 -7195
rect 7687 -7256 7692 -7200
rect 7748 -7256 7753 -7200
rect 7687 -7261 7753 -7256
rect 8362 -7486 8478 -7481
rect 8362 -7582 8372 -7486
rect 8468 -7582 8478 -7486
rect 8362 -7587 8478 -7582
<< via3 >>
rect 5042 984 5138 1080
rect 5062 -256 5158 -160
rect 5032 -1056 5128 -960
rect 5052 -1856 5148 -1760
rect 5046 -2655 5142 -2559
rect 5062 -3456 5158 -3360
rect 5036 -4256 5132 -4160
rect 5036 -5056 5132 -4960
rect 5032 -5856 5128 -5760
rect 5032 -7044 5128 -6948
rect 8416 440 8512 536
rect 8386 -800 8482 -704
rect 8398 -1600 8494 -1504
rect 8396 -2400 8492 -2304
rect 8380 -3200 8476 -3104
rect 8370 -4000 8466 -3904
rect 8388 -4800 8484 -4704
rect 8370 -5600 8466 -5504
rect 8394 -6399 8490 -6303
rect 8372 -7582 8468 -7486
<< metal4 >>
rect 4854 1080 5322 1266
rect 4854 984 5042 1080
rect 5138 984 5322 1080
rect 4854 -160 5322 984
rect 4854 -256 5062 -160
rect 5158 -256 5322 -160
rect 4854 -960 5322 -256
rect 4854 -1056 5032 -960
rect 5128 -1056 5322 -960
rect 4854 -1760 5322 -1056
rect 4854 -1856 5052 -1760
rect 5148 -1856 5322 -1760
rect 4854 -2559 5322 -1856
rect 4854 -2655 5046 -2559
rect 5142 -2655 5322 -2559
rect 4854 -3360 5322 -2655
rect 4854 -3456 5062 -3360
rect 5158 -3456 5322 -3360
rect 4854 -4160 5322 -3456
rect 4854 -4256 5036 -4160
rect 5132 -4256 5322 -4160
rect 4854 -4960 5322 -4256
rect 4854 -5056 5036 -4960
rect 5132 -5056 5322 -4960
rect 4854 -5760 5322 -5056
rect 4854 -5856 5032 -5760
rect 5128 -5856 5322 -5760
rect 4854 -6948 5322 -5856
rect 4854 -7044 5032 -6948
rect 5128 -7044 5322 -6948
rect 4854 -7118 5322 -7044
rect 8186 536 8654 738
rect 8186 440 8416 536
rect 8512 440 8654 536
rect 8186 -704 8654 440
rect 8186 -800 8386 -704
rect 8482 -800 8654 -704
rect 8186 -1504 8654 -800
rect 8186 -1600 8398 -1504
rect 8494 -1600 8654 -1504
rect 8186 -2304 8654 -1600
rect 8186 -2400 8396 -2304
rect 8492 -2400 8654 -2304
rect 8186 -3104 8654 -2400
rect 8186 -3200 8380 -3104
rect 8476 -3200 8654 -3104
rect 8186 -3904 8654 -3200
rect 8186 -4000 8370 -3904
rect 8466 -4000 8654 -3904
rect 8186 -4704 8654 -4000
rect 8186 -4800 8388 -4704
rect 8484 -4800 8654 -4704
rect 8186 -5504 8654 -4800
rect 8186 -5600 8370 -5504
rect 8466 -5600 8654 -5504
rect 8186 -6303 8654 -5600
rect 8186 -6399 8394 -6303
rect 8490 -6399 8654 -6303
rect 8186 -7486 8654 -6399
rect 8186 -7582 8372 -7486
rect 8468 -7582 8654 -7486
rect 8186 -7646 8654 -7582
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683272759
transform 1 0 5438 0 1 -3152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1683272759
transform 1 0 5438 0 1 -6352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1683272759
transform 1 0 5438 0 1 -1552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1683272759
transform 1 0 5438 0 1 -2352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1683272759
transform 1 0 5438 0 1 -752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1683272759
transform 1 0 5438 0 1 -3952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1683272759
transform 1 0 5438 0 1 -4752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1683272759
transform 1 0 7782 0 1 -6352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1683272759
transform 1 0 7782 0 1 -5552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_9
timestamp 1683272759
transform 1 0 7782 0 1 -4752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_10
timestamp 1683272759
transform 1 0 7782 0 1 -3952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_11
timestamp 1683272759
transform 1 0 7782 0 1 -3152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_12
timestamp 1683272759
transform 1 0 7782 0 1 -2352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_13
timestamp 1683272759
transform 1 0 7782 0 1 -1552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_14
timestamp 1683272759
transform 1 0 7782 0 1 -752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_15
timestamp 1683272759
transform 1 0 5438 0 1 -5552
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  x1
timestamp 1683272759
transform 1 0 5790 0 1 -752
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x2
timestamp 1683272759
transform 1 0 5790 0 1 -1552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x3
timestamp 1683272759
transform 1 0 5790 0 1 -2352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x4
timestamp 1683272759
transform 1 0 5790 0 1 -3152
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x5
timestamp 1683272759
transform 1 0 5790 0 1 -3952
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x6
timestamp 1683272759
transform 1 0 5790 0 1 -4752
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x7
timestamp 1683272759
transform 1 0 5790 0 1 -5552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x8
timestamp 1683272759
transform 1 0 5790 0 1 -6352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x9
timestamp 1683272759
transform 1 0 6786 0 1 -6352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x10
timestamp 1683272759
transform 1 0 6786 0 1 -5552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x11
timestamp 1683272759
transform 1 0 6786 0 1 -4752
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x12
timestamp 1683272759
transform 1 0 6786 0 1 -3952
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x13
timestamp 1683272759
transform 1 0 6786 0 1 -3152
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x14
timestamp 1683272759
transform 1 0 6786 0 1 -2352
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x15
timestamp 1683272759
transform 1 0 6786 0 1 -1552
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_2  x16
timestamp 1683272759
transform 1 0 6786 0 1 -752
box -38 -48 958 592
use sky130_fd_sc_hd__inv_8  x17 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683272759
transform 1 0 6785 0 1 -7533
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x18
timestamp 1683272759
transform 1 0 5881 0 1 -7533
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x19
timestamp 1683272759
transform 1 0 6762 0 1 488
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x20
timestamp 1683272759
transform 1 0 5858 0 1 488
box -38 -48 866 592
<< labels >>
rlabel metal3 6000 240 6060 300 1 S1
port 2 n
rlabel metal3 6130 240 6190 300 1 S1N
rlabel metal3 6260 240 6320 300 1 S2
port 1 n
rlabel metal3 6390 240 6450 300 1 S2N
rlabel metal3 6520 240 6580 300 1 S3
port 0 n
rlabel metal3 6650 240 6710 300 1 S3N
rlabel metal3 5870 240 5930 300 1 S0N
rlabel metal3 5740 240 5800 300 1 S0
port 39 n
flabel metal1 7700 968 7900 1168 0 FreeSans 256 0 0 0 VPWR
port 5 nsew
flabel metal1 5606 -7634 5806 -7434 0 FreeSans 256 0 0 0 VGND
port 4 nsew
flabel metal1 4338 -776 4538 -576 0 FreeSans 256 180 0 0 Q0
port 37 nsew
flabel metal1 4334 -520 4534 -320 0 FreeSans 256 0 0 0 Q0N
port 21 nsew
flabel metal1 4372 -1248 4572 -1048 0 FreeSans 256 0 0 0 Q1N
port 20 nsew
flabel metal1 4314 -2070 4514 -1870 0 FreeSans 256 0 0 0 Q2N
port 18 nsew
flabel metal1 4336 -2876 4536 -2676 0 FreeSans 256 0 0 0 Q3N
port 17 nsew
flabel metal1 4356 -3636 4556 -3436 0 FreeSans 256 0 0 0 Q4N
port 16 nsew
flabel metal1 4348 -4460 4548 -4260 0 FreeSans 256 0 0 0 Q5N
port 22 nsew
flabel metal1 4350 -5310 4550 -5110 0 FreeSans 256 0 0 0 Q6N
port 15 nsew
flabel metal1 4324 -6036 4524 -5836 0 FreeSans 256 0 0 0 Q7N
port 14 nsew
flabel metal1 4376 -1546 4576 -1346 0 FreeSans 256 180 0 0 Q1
port 36 nsew
flabel metal1 4376 -2324 4576 -2124 0 FreeSans 256 180 0 0 Q2
port 35 nsew
flabel metal1 4366 -3148 4566 -2948 0 FreeSans 256 180 0 0 Q3
port 34 nsew
flabel metal1 4366 -3896 4566 -3696 0 FreeSans 256 180 0 0 Q4
port 33 nsew
flabel metal1 4386 -4752 4586 -4552 0 FreeSans 256 0 0 0 Q5
port 38 nsew
flabel metal1 4356 -5558 4556 -5358 0 FreeSans 256 180 0 0 Q6
port 32 nsew
flabel metal1 4366 -6324 4566 -6124 0 FreeSans 256 180 0 0 Q7
port 31 nsew
flabel metal1 9354 -6048 9554 -5848 0 FreeSans 256 0 0 0 Q8N
port 13 nsew
flabel metal1 9374 -5235 9574 -5035 0 FreeSans 256 0 0 0 Q9N
port 12 nsew
flabel metal1 9352 -2873 9552 -2673 0 FreeSans 256 0 0 0 Q12N
port 9 nsew
flabel metal1 9320 -2092 9520 -1892 0 FreeSans 256 0 0 0 Q13N
port 8 nsew
flabel metal1 9206 -1280 9406 -1080 0 FreeSans 256 0 0 0 Q14N
port 6 nsew
flabel metal1 9310 -484 9510 -284 0 FreeSans 256 0 0 0 Q15N
port 7 nsew
flabel metal1 9320 -3654 9520 -3454 0 FreeSans 256 0 0 0 Q11N
port 11 nsew
flabel metal1 9246 -4470 9446 -4270 0 FreeSans 256 0 0 0 Q10N
port 10 nsew
flabel metal1 8842 -3082 9042 -2882 0 FreeSans 256 0 0 0 Q12
port 26 nsew
flabel metal1 8814 -2268 9014 -2068 0 FreeSans 256 0 0 0 Q13
port 25 nsew
flabel metal1 8754 -1472 8954 -1272 0 FreeSans 256 0 0 0 Q14
port 23 nsew
flabel metal1 8732 -660 8932 -460 0 FreeSans 256 0 0 0 Q15
port 24 nsew
flabel metal1 8878 -4666 9078 -4466 0 FreeSans 256 0 0 0 Q10
port 27 nsew
flabel metal1 8862 -3864 9062 -3664 0 FreeSans 256 0 0 0 Q11
port 28 nsew
flabel metal1 8892 -6260 9092 -6060 0 FreeSans 256 0 0 0 Q8
port 30 nsew
flabel metal1 8942 -5466 9142 -5266 0 FreeSans 256 0 0 0 Q9
port 29 nsew
<< end >>
