** sch_path: /foss/designs/analog_mux_files/decoder_x4.sch

.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt decoder_x4 S3 S2 S1 S0 VGND VPWR Q14N Q15N Q13N Q12N Q10N Q11N Q9N Q8N Q7N Q6N Q4N Q3N Q2N
+ Q1N Q0N Q5N Q14 Q15 Q13 Q12 Q10 Q11 Q9 Q8 Q7 Q6 Q4 Q3 Q2 Q1 Q0 Q5
*.PININFO S3:I S2:I S1:I S0:I VGND:I VPWR:I Q14N:O Q15N:O Q13N:O Q12N:O Q10N:O Q11N:O Q9N:O Q8N:O
*+ Q7N:O Q6N:O Q4N:O Q3N:O Q2N:O Q1N:O Q0N:O Q5N:O Q14:O Q15:O Q13:O Q12:O Q10:O Q11:O Q9:O Q8:O Q7:O Q6:O
*+ Q4:O Q3:O Q2:O Q1:O Q0:O Q5:O
x17 S3 VGND VGND VPWR VPWR S3N sky130_fd_sc_hd__inv_8
x18 S2 VGND VGND VPWR VPWR S2N sky130_fd_sc_hd__inv_8
x19 S1 VGND VGND VPWR VPWR S1N sky130_fd_sc_hd__inv_8
x20 S0 VGND VGND VPWR VPWR S0N sky130_fd_sc_hd__inv_8
x21 Q0N VGND VGND VPWR VPWR Q0 sky130_fd_sc_hd__inv_2
x22 Q1N VGND VGND VPWR VPWR Q1 sky130_fd_sc_hd__inv_2
x23 Q2N VGND VGND VPWR VPWR Q2 sky130_fd_sc_hd__inv_2
x24 Q3N VGND VGND VPWR VPWR Q3 sky130_fd_sc_hd__inv_2
x1 S3N S2N S1N S0N VGND VGND VPWR VPWR Q0N sky130_fd_sc_hd__nand4_2
x2 S3N S2N S1N S0 VGND VGND VPWR VPWR Q1N sky130_fd_sc_hd__nand4_2
x3 S3N S2N S1 S0N VGND VGND VPWR VPWR Q2N sky130_fd_sc_hd__nand4_2
x4 S3N S2N S1 S0 VGND VGND VPWR VPWR Q3N sky130_fd_sc_hd__nand4_2
x5 S3N S2 S1N S0N VGND VGND VPWR VPWR Q4N sky130_fd_sc_hd__nand4_2
x6 S3N S2 S1N S0 VGND VGND VPWR VPWR Q5N sky130_fd_sc_hd__nand4_2
x7 S3N S2 S1 S0N VGND VGND VPWR VPWR Q6N sky130_fd_sc_hd__nand4_2
x8 S3N S2 S1 S0 VGND VGND VPWR VPWR Q7N sky130_fd_sc_hd__nand4_2
x9 S3 S2N S1N S0N VGND VGND VPWR VPWR Q8N sky130_fd_sc_hd__nand4_2
x10 S3 S2N S1N S0 VGND VGND VPWR VPWR Q9N sky130_fd_sc_hd__nand4_2
x11 S3 S2N S1 S0N VGND VGND VPWR VPWR Q10N sky130_fd_sc_hd__nand4_2
x12 S3 S2N S1 S0 VGND VGND VPWR VPWR Q11N sky130_fd_sc_hd__nand4_2
x13 S3 S2 S1N S0N VGND VGND VPWR VPWR Q12N sky130_fd_sc_hd__nand4_2
x14 S3 S2 S1N S0 VGND VGND VPWR VPWR Q13N sky130_fd_sc_hd__nand4_2
x15 S3 S2 S1 S0N VGND VGND VPWR VPWR Q14N sky130_fd_sc_hd__nand4_2
x16 S3 S2 S1 S0 VGND VGND VPWR VPWR Q15N sky130_fd_sc_hd__nand4_2
x25 Q4N VGND VGND VPWR VPWR Q4 sky130_fd_sc_hd__inv_2
x26 Q5N VGND VGND VPWR VPWR Q5 sky130_fd_sc_hd__inv_2
x27 Q6N VGND VGND VPWR VPWR Q6 sky130_fd_sc_hd__inv_2
x28 Q7N VGND VGND VPWR VPWR Q7 sky130_fd_sc_hd__inv_2
x29 Q8N VGND VGND VPWR VPWR Q8 sky130_fd_sc_hd__inv_2
x30 Q9N VGND VGND VPWR VPWR Q9 sky130_fd_sc_hd__inv_2
x31 Q10N VGND VGND VPWR VPWR Q10 sky130_fd_sc_hd__inv_2
x32 Q11N VGND VGND VPWR VPWR Q11 sky130_fd_sc_hd__inv_2
x33 Q12N VGND VGND VPWR VPWR Q12 sky130_fd_sc_hd__inv_2
x34 Q13N VGND VGND VPWR VPWR Q13 sky130_fd_sc_hd__inv_2
x35 Q14N VGND VGND VPWR VPWR Q14 sky130_fd_sc_hd__inv_2
x36 Q15N VGND VGND VPWR VPWR Q15 sky130_fd_sc_hd__inv_2
.ends
.end
