* NGSPICE file created from decoder_x4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VPWR Y VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=2.05e+12p pd=1.41e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=5.915e+11p pd=5.72e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt decoder_x4 S3 S2 S1 VGND VPWR Q14N Q15N Q13N Q12N Q10N Q11N Q9N Q8N Q7N Q6N
+ Q4N Q3N Q2N Q1N Q0N Q5N Q14 Q15 Q13 Q12 Q10 Q11 Q9 Q8 Q7 Q6 Q4 Q3 Q2 Q1 Q0 Q5 S0
Xx1 S3N S2N S1N S0N VGND VPWR Q0N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx2 S3N S2N S1N S0 VGND VPWR Q1N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx3 S3N S2N S1 S0N VGND VPWR Q2N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx4 S3N S2N S1 S0 VGND VPWR Q3N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx5 S3N S2 S1N S0N VGND VPWR Q4N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx6 S3N S2 S1N S0 VGND VPWR Q5N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx7 S3N S2 S1 S0N VGND VPWR Q6N VGND VPWR sky130_fd_sc_hd__nand4_2
Xsky130_fd_sc_hd__inv_2_11 Q12N VGND VPWR Q12 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_10 Q11N VGND VPWR Q11 VGND VPWR sky130_fd_sc_hd__inv_2
Xx8 S3N S2 S1 S0 VGND VPWR Q7N VGND VPWR sky130_fd_sc_hd__nand4_2
Xsky130_fd_sc_hd__inv_2_12 Q13N VGND VPWR Q13 VGND VPWR sky130_fd_sc_hd__inv_2
Xx9 S3 S2N S1N S0N VGND VPWR Q8N VGND VPWR sky130_fd_sc_hd__nand4_2
Xsky130_fd_sc_hd__inv_2_13 Q14N VGND VPWR Q14 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_14 Q15N VGND VPWR Q15 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_0 Q3N VGND VPWR Q3 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_15 Q6N VGND VPWR Q6 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 Q7N VGND VPWR Q7 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_2 Q1N VGND VPWR Q1 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_3 Q2N VGND VPWR Q2 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_4 Q0N VGND VPWR Q0 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_5 Q4N VGND VPWR Q4 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_6 Q5N VGND VPWR Q5 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_7 Q8N VGND VPWR Q8 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_8 Q9N VGND VPWR Q9 VGND VPWR sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_9 Q10N VGND VPWR Q10 VGND VPWR sky130_fd_sc_hd__inv_2
Xx20 S0 VGND VPWR S0N VGND VPWR sky130_fd_sc_hd__inv_8
Xx10 S3 S2N S1N S0 VGND VPWR Q9N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx11 S3 S2N S1 S0N VGND VPWR Q10N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx12 S3 S2N S1 S0 VGND VPWR Q11N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx13 S3 S2 S1N S0N VGND VPWR Q12N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx15 S3 S2 S1 S0N VGND VPWR Q14N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx14 S3 S2 S1N S0 VGND VPWR Q13N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx16 S3 S2 S1 S0 VGND VPWR Q15N VGND VPWR sky130_fd_sc_hd__nand4_2
Xx17 S3 VGND VPWR S3N VGND VPWR sky130_fd_sc_hd__inv_8
Xx18 S2 VGND VPWR S2N VGND VPWR sky130_fd_sc_hd__inv_8
Xx19 S1 VGND VPWR S1N VGND VPWR sky130_fd_sc_hd__inv_8
.ends

